`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/10/24 16:59:56
// Design Name: 
// Module Name: reg8file
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module reg8file (
    input  wire clk,  
    input  wire clr,    
    input  wire en,
    input  wire [7:0] d,
    input  wire [2:0] wsel,
    input  wire [2:0] rsel,
    output reg  [7:0] q    
);
reg [7:0] regfile [7:0];
always @(posedge clk or posedge clr) begin
    if (clr == 1'b1) begin
        // ��λʱ������8���Ĵ���ֱ�����㣨����ʱ�ӣ��첽��Ч��
        regfile[0] <= 8'b0;
        regfile[1] <= 8'b0;
        regfile[2] <= 8'b0;
        regfile[3] <= 8'b0;
        regfile[4] <= 8'b0;
        regfile[5] <= 8'b0;
        regfile[6] <= 8'b0;
        regfile[7] <= 8'b0;
    end else if (en == 1'b1) begin
        // дʹ����Чʱ����ʱ�������أ�������dд��wselָ���ļĴ���
        regfile[wsel] <= d;
    end
    // ��en=0����ִ��д�������Ĵ�������ԭ��ֵ�����������룬Ĭ����Ϊ��
end

// ����߼����첽����������ַ�仯ʱ������������£�
always @(*) begin
    q = regfile[rsel]; // ֱ�Ӷ�ȡrselָ���ļĴ���ֵ����ʱ���ӳ�
end

endmodule
