`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/10/24 16:00:13
// Design Name: 
// Module Name: dff
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module dff (
    input      clk,
    input      clr,
    input      en ,
    input      d  ,
    output reg q
);
always @(posedge clk or posedge clr) begin
    if (clr == 1'b1) begin  // ��һ�����ȿ������ź��Ƿ���Ч��1'b1��ʾ������1��
        q <= 1'b0;          // ���㣺qֱ�ӱ��0��<=��ʱ��ֵ�������������
    end
    else if (en == 1'b1) begin  // �ڶ�������������㣬��ʹ���Ƿ�����
        q <= d;                 // ������ʱ�������أ���d��ֵ����q�������ݣ�
    end
end
endmodule
