`timescale 1ns / 1ps

module uart_recv(
    input clk,
    input rst,
    input din,
    output reg valid,
    output reg [7:0] data
);

    // ״̬����
    localparam IDLE  = 3'b000;
    localparam START = 3'b001;
    localparam DATA  = 3'b010;
    localparam STOP  = 3'b011;
    
    // �����ʲ��� - ��������
    localparam CLK_FREQ = 100_000_000;//100MHz
    localparam BAUD_RATE = 9600;//������
    localparam BIT_CYCLES = CLK_FREQ / BAUD_RATE;  // 10416
    localparam BIT_CYCLES_HALF = BIT_CYCLES / 2;   // 5208
    
    // ״̬�Ĵ���
    reg [2:0] current_state, next_state;
    
    // ������
    reg [13:0] bit_counter;
    reg [2:0] bit_index;
    reg [7:0] data_shift;
    
    // ����ͬ���Ĵ�������ֹ����̬
     reg din_sync1, din_sync2, din_sync3;
    
      always @(posedge clk or posedge rst) begin
        if (rst) begin
            din_sync1 <= 1'b1;
            din_sync2 <= 1'b1;
            din_sync3 <= 1'b1;
        end else begin
            din_sync1 <= din;      // ��һ��ͬ��
            din_sync2 <= din_sync1; // �ڶ���ͬ��
            din_sync3 <= din_sync2; // ������ͬ��
        end
    end
    
    // ==================== ״̬ת���߼� ====================
    always @(posedge clk or posedge rst) begin
        if (rst) 
            current_state <= IDLE;
        else 
            current_state <= next_state;
    end
    
    // ==================== ��һ״̬�߼� ====================
    always @(*) begin
        case (current_state)
            IDLE:  next_state = (!din_sync2) ? START : IDLE;  // �����ʼλ
            START: next_state = (bit_counter == BIT_CYCLES - 1) ? DATA : START;  // ��������
            DATA:  next_state = (bit_index == 3'd7 && bit_counter == BIT_CYCLES - 1) ? STOP : DATA;
            STOP:  next_state = (bit_counter == BIT_CYCLES - 1) ? IDLE : STOP;
            default: next_state = IDLE;
        endcase
    end
    
    // ==================== λ���������� ====================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            bit_counter <= 0;
        end else begin
            case (current_state)
                IDLE: begin
                    bit_counter <= 0;
                end
                
                START, DATA, STOP: begin
                    if (bit_counter < BIT_CYCLES - 1)
                        bit_counter <= bit_counter + 1;
                    else
                        bit_counter <= 0;
                end
                
                default: begin
                    bit_counter <= 0;
                end
            endcase
        end
    end
    
    // ==================== λ�������� ====================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            bit_index <= 0;
        end else begin
            if (current_state == DATA) begin
                if (bit_counter == BIT_CYCLES - 1) begin
                    if (bit_index < 3'd7)
                        bit_index <= bit_index + 1;
                    else
                        bit_index <= 0;
                end
            end else begin
                bit_index <= 0;
            end
        end
    end
    
    // ==================== ������λ���� ====================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            data_shift <= 0;
        end else begin
            if (current_state == DATA) begin
                if (bit_counter == BIT_CYCLES_HALF - 1) begin  // ������λ�м����
                    data_shift <= {din_sync3, data_shift[7:1]};
                end
            end else if (current_state == IDLE) begin
                data_shift <= 0;
            end
        end
    end
   
    // ==================== ��Ч�źſ��� ====================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            valid <= 1'b0;
        end else begin
            valid <= 1'b0;  // Ĭ��validΪ0
            
            if (current_state == STOP) begin
                if (bit_counter == BIT_CYCLES_HALF - 1) begin
                    valid <= 1'b1;  // ��ֹͣλ�м�ʱ�������Ч����
                end
            end
        end
    end
    
    // ==================== ����������� ====================
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            data <= 8'b0;
        end else begin
            if (current_state == STOP) begin
                if (bit_counter == BIT_CYCLES_HALF - 1) begin
                    data <= data_shift;  // ��ֹͣλ�м�ʱ���������
                end
            end
        end
    end

endmodule