`timescale 1ns / 1ps

module reg8file_tb ();

    reg clk;
    reg clr;
    reg en;
    reg [2:0] wsel;  
    reg [2:0] rsel;  
    reg [7:0] d;
    wire [7:0] q;

    reg8file u_reg8file (
        .clk(clk),   // ʱ������
        .clr(clr),   // ��λ����
        .en(en),     // дʹ������
        .wsel(wsel), // д��ַ����
        .rsel(rsel), // ����ַ����
        .d(d),       // д����������
        .q(q)        // ������������
    );


    initial begin
        clk = 1'b0;          // ��ʼʱ��Ϊ0
        forever #10 clk = ~clk; // ÿ10ns��תһ�Σ�ʱ������20ns��50MHz��
    end

    // ------------------- ���Լ������� -------------------
    initial begin
        // �׶�1����λ���ԣ��첽�������мĴ�����
        clr = 1'b1;  // ��λ��Ч���ߵ�ƽ��
        en  = 1'b0;  // дʹ�ܹر�
        wsel = 3'b000;
        rsel = 3'b000;
        d    = 8'h00;
        #20;  // �ȴ�20ns��1��ʱ�����ڣ����۲츴λЧ��

        // �׶�2��д�������ԣ���ͬ�Ĵ���д�����ݣ�
        clr = 1'b0;  // �ͷŸ�λ
        en  = 1'b1;  // ʹ��д����

        wsel = 3'b000; // д����0�żĴ�����
        d    = 8'hAA;  // д������0xAA
        #20;           // ʱ�������ش���д����

        wsel = 3'b001; // д����1�żĴ�����
        d    = 8'h55;  // д������0x55
        #20;

        wsel = 3'b010; // д����2�żĴ�����
        d    = 8'hFF;  // д������0xFF
        #20;

        // �׶�3�����������ԣ��ر�дʹ�ܣ�����ͬ�Ĵ�����
        en = 1'b0;     // �ر�дʹ��

        rsel = 3'b000; // ������0�żĴ�������Ԥ��q=0xAA��
        #20;

        rsel = 3'b001; // ������1�żĴ�������Ԥ��q=0x55��
        #20;

        rsel = 3'b010; // ������2�żĴ�������Ԥ��q=0xFF��
        #20;

        // �׶�4������д���ԣ�����д��0�żĴ�����
        en = 1'b1;
        wsel = 3'b000;
        d    = 8'hCC;  // д��������0xCC
        #20;

        en = 1'b0;
        rsel = 3'b000; // ������0�żĴ�������Ԥ��q=0xCC��
        #20;

        // �׶�5���ٴθ�λ���ԣ���֤�첽���㣩
        clr = 1'b1;    // ��λ��Ч
        #20;

        clr = 1'b0;
        rsel = 3'b000; // ������0�żĴ�������Ԥ��q=0x00��
        #20;

        $finish; // ��������
    end

    // ------------------- ���Ը�������ӡ�ź� -------------------
    always @(posedge clk) begin
        $display("Time=%t: clr=%b, en=%b, wsel=%b, rsel=%b, d=%h, q=%h", 
                 $time, clr, en, wsel, rsel, d, q);
    end

endmodule