
module top(
    input wire clk,
    input wire sw0,
    input wire s1,     // S1��Ϊ�첽��λ
    input wire s2,     // S2��Ϊ��������ͣ����
    input wire s3,     // S3��Ϊ��������
    output wire [7:0] led_en,
    output wire [7:0] led_cx
);

    // ѧ�ź���λ
    localparam STUDENT_ID_HIGH = 4'h6;  // ѧ��ʮλ
    localparam STUDENT_ID_LOW  = 4'h8;  // ѧ�Ÿ�λ

    // �ڲ��źŶ���
    wire [6:0] count_no_debounce;    // ���������� (0-99)
    wire [6:0] count_with_debounce;  // ���������� (0-99)
    wire [4:0] decimal_count;        // ʮ���Ƽ��� (0-30)
    wire [3:0] decimal_ten;          // ʮ����ʮλ
    wire [3:0] decimal_unit;         // ʮ���Ƹ�λ
    wire debounced_s3;               // �������S3�ź�
    wire debounced_s2;               // �������S2�ź�
    wire s3_edge;                    // S3���ؼ��
    wire s3_debounced_edge;          // ������S3���ؼ��
    wire s2_debounced_edge;          // ������S2���ؼ��
    wire counter_enable;             // ������ʹ��
    
    // S2��������ģ��ʵ����
    debounce u_debounce_s2(
        .clk(clk),
        .rst(s1),
        .key_in(s2),
        .key_out(debounced_s2)
    );
    
    // S3��������ģ��ʵ����
    debounce u_debounce_s3(
        .clk(clk),
        .rst(s1),
        .key_in(s3),
        .key_out(debounced_s3)
    );
    
    // ���ؼ��ģ��ʵ����
    edge_detector u_edge_detector_s3(
        .clk(clk),
        .rst(s1),
        .signal_in(s3),
        .pos_edge(s3_edge)
    );
    
    edge_detector u_edge_detector_s3_debounced(
        .clk(clk),
        .rst(s1),
        .signal_in(debounced_s3),
        .pos_edge(s3_debounced_edge)
    );
    
    edge_detector u_edge_detector_s2_debounced(
        .clk(clk),
        .rst(s1),
        .signal_in(debounced_s2),
        .pos_edge(s2_debounced_edge)
    );
    
    // ������������ (0-99)
    counter_0to99 u_counter_no_debounce(
        .clk(clk),
        .rst(s1),
        .en(s3_edge),           // ʹ��δ�����ı����ź�
        .count(count_no_debounce)
    );
    
    // ������������ (0-99)
    counter_0to99 u_counter_with_debounce(
        .clk(clk),
        .rst(s1),
        .en(s3_debounced_edge), // ʹ��������ı����ź�
        .count(count_with_debounce)
    );
    
    // ʮ���Ƽ���������
    toggle_ff u_toggle_ff(
        .clk(clk),
        .rst(s1),
        .toggle(s2_debounced_edge),
        .out(counter_enable)
    );
    
    // 0.1s�����0-30������
    decimal_counter u_decimal_counter(
        .clk(clk),
        .rst(s1),
        .enable(counter_enable),
        .count(decimal_count),
        .display_ten(decimal_ten),
        .display_unit(decimal_unit)
    );
    
    // ��7λ���������Ϊʮλ�͸�λ��ʾ (0-99)
    wire [3:0] no_debounce_ten;   // ����������ʮλ
    wire [3:0] no_debounce_unit;  // ������������λ
    wire [3:0] with_debounce_ten; // ����������ʮλ  
    wire [3:0] with_debounce_unit;// ������������λ
    
    // 7λ������ֵ���Ϊʮλ�͸�λ (0-99)
    assign no_debounce_ten = count_no_debounce / 7'd10;
    assign no_debounce_unit = count_no_debounce % 7'd10;
    
    assign with_debounce_ten = count_with_debounce / 7'd10;
    assign with_debounce_unit = count_with_debounce % 7'd10;
    
    // �������ʾ�������
    wire [31:0] display_data;
    assign display_data = {
        STUDENT_ID_HIGH,        // DK7 - ѧ��ʮλ
        STUDENT_ID_LOW,         // DK6 - ѧ�Ÿ�λ
        no_debounce_ten,        // DK5 - ����������ʮλ
        no_debounce_unit,       // DK4 - ������������λ
        with_debounce_ten,      // DK3 - ����������ʮλ
        with_debounce_unit,     // DK2 - ������������λ
        decimal_ten,            // DK1 - ʮ���Ƽ���ʮλ
        decimal_unit            // DK0 - ʮ���Ƽ�����λ
    };
    
    // ����ܿ���ģ��
    led_ctrl_unit u_led_ctrl_unit(
        .rst(s1),
        .clk(clk),
        .display(display_data),
        .enable(sw0),
        .led_en(led_en),
        .led_cx(led_cx)
    );

endmodule
